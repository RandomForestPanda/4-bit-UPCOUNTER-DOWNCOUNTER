module and(
    
);
    
endmodule